`timescale 1ps / 1ps
module test_Code_generation;

wire [15:0] D_out;
reg [28:0] INST;
wire Over_Flow;
ALU alu(INST,D_out,Over_Flow);

initial	// Test stimulus
  begin
    #0   INST = 29'b00101000100000000000000000000; //addi $R1, $R0, 0 
		#350 INST = 29'b00101001000000000000000000000; //addi $R2, $R0, 0

		#350 INST = 29'b00100000100010010000000000000; //add $R1, $R1, $R2
		#350 INST = 29'b00101001000100000000000000001; //addi $R2, $R2, 1

		#350 INST = 29'b00100000100010010000000000000; //add $R1, $R1, $R2
		#350 INST = 29'b00101001000100000000000000001; //addi $R2, $R2, 1

		#350 INST = 29'b00100000100010010000000000000; //add $R1, $R1, $R2
		#350 INST = 29'b00101001000100000000000000001; //addi $R2, $R2, 1

		#350 INST = 29'b00100000100010010000000000000; //add $R1, $R1, $R2
		#350 INST = 29'b00101001000100000000000000001; //addi $R2, $R2, 1

		#350 INST = 29'b00100000100010010000000000000; //add $R1, $R1, $R2
		#350 INST = 29'b00101001000100000000000000001; //addi $R2, $R2, 1

		#350 INST = 29'b00100000100010010000000000000; //add $R1, $R1, $R2
		#350 INST = 29'b00101001000100000000000000001; //addi $R2, $R2, 1

		#350 INST = 29'b00100000100010010000000000000; //add $R1, $R1, $R2
		#350 INST = 29'b00101001000100000000000000001; //addi $R2, $R2, 1

		#350 INST = 29'b00100000100010010000000000000; //add $R1, $R1, $R2
		#350 INST = 29'b00101001000100000000000000001; //addi $R2, $R2, 1

		#350 INST = 29'b00100000100010010000000000000; //add $R1, $R1, $R2
		#350 INST = 29'b00101001000100000000000000001; //addi $R2, $R2, 1

		#350 INST = 29'b00100000100010010000000000000; //add $R1, $R1, $R2
		#350 INST = 29'b00101001000100000000000000001; //addi $R2, $R2, 1
 
  end

endmodule 